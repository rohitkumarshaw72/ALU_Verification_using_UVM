
package alu_pkg;

    import uvm_pkg::*;
    
    `include "uvm_macros.svh"
    
    `include "alu_xtn.sv"
    `include "alu_config.sv"
    `include "env_config.sv"
    
    `include "alu_driver.sv"
    `include "alu_monitor.sv"
    `include "alu_seqr.sv"
    `include "alu_write_agent.sv"
    `include "alu_write_agent_top.sv"
    `include "alu_seq.sv"
    
    `include "alu_virtual_seqr.sv"
    `include "alu_virtual_seq.sv"
    `include "alu_scoreboard.sv"
    
    `include "alu_env.sv"
    
    `include "alu_test.sv"

endpackage
